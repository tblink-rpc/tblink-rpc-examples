/****************************************************************************
 * py_uvm_seq_tb.sv
 ****************************************************************************/

  
/**
 * Module: py_uvm_seq_tb
 * 
 * TODO: Add module documentation
 */
module py_uvm_seq_tb;
	import uvm_pkg::*;
	import py_uvm_seq_pkg::*;
	
	initial begin
		run_test();
	end

endmodule


