/****************************************************************************
 * my_seq_2.svh
 ****************************************************************************/

  
/**
 * Class: my_seq_2
 * 
 * TODO: Add class documentation
 */
class my_seq_2 extends my_seq_2_if_base #(my_seq_base);

	function new(string name="my_seq_2");
		super.new(name);
	endfunction


endclass


