
/****************************************************************************
 * my_seq_1.svh
 ****************************************************************************/

  
/**
 * Class: my_seq_1
 * 
 * TODO: Add class documentation
 */
class my_seq_1 extends my_seq_1_if_base #(my_seq_base);
	`uvm_object_utils(my_seq_1)

	function new(string name="py_uvm_seq");
		super.new(name);
	endfunction


endclass


