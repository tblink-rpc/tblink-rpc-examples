/****************************************************************************
 * py_uvm_seq_pkg.sv
 ****************************************************************************/
`include "uvm_macros.svh"
  
/**
 * Package: py_uvm_seq_pkg
 * 
 * TODO: Add package documentation
 */
package py_uvm_seq_pkg;
	import uvm_pkg::*;
	import tblink_rpc_uvm::*;

	`include "my_seq_if.svh"
	`include "py_uvm_seq.svh"
	`include "py_uvm_seq_test.svh"

endpackage


